//-------------------------------------------------------------------------
//						fpu_agent - www.verificationguide.com 
//-------------------------------------------------------------------------

`include "fpu_seq_item.sv"
`include "fpu_sequencer.sv"
`include "fpu_sequence.sv"
`include "fpu_driver.sv"
`include "fpu_monitor.sv"

class fpu_agent extends uvm_agent;

  //---------------------------------------
  // component instances
  //---------------------------------------
  fpu_driver    driver;
  fpu_sequencer sequencer;
  fpu_monitor   monitor;

  `uvm_component_utils(fpu_agent)
  
  //---------------------------------------
  // constructor
  //---------------------------------------
  function new (string name, uvm_component parent);
    super.new(name, parent);
  endfunction : new

  //---------------------------------------
  // build_phase
  //---------------------------------------
  function void build_phase(uvm_phase phase);
    super.build_phase(phase);
    
    monitor = fpu_monitor::type_id::create("monitor", this);

    //creating driver and sequencer only for ACTIVE agent
    if(get_is_active() == UVM_ACTIVE) begin
      driver    = fpu_driver::type_id::create("driver", this);
      sequencer = fpu_sequencer::type_id::create("sequencer", this);
    end
  endfunction : build_phase
  
  //---------------------------------------  
  // connect_phase - connecting the driver and sequencer port
  //---------------------------------------
  function void connect_phase(uvm_phase phase);
    if(get_is_active() == UVM_ACTIVE) begin
      driver.seq_item_port.connect(sequencer.seq_item_export);
    end
  endfunction : connect_phase

endclass : fpu_agent