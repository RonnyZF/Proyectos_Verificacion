`include "interface.sv"
`include "stimulus.sv"
`include "scoreboard.sv"
`include "driver.sv"
`include "monitor.sv"
`include "env.sv"
`include "test_1.sv"
`include "assertions.sv"
//`include "test_2.sv"
`include "top.sv"
