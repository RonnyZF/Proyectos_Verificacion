`include "except.v"
`include "post_norm.v"
`include "pre_norm.v"
`include "pre_norm_fmul.v"
`include "primitives.v"
`include "fpu.v"
