class scoreboard;
  logic [7:0] store [$];
endclass
