
class scoreboard;
  logic [31:0] opa [$];
  logic [31:0] opb [$];
endclass
